`timescale 1 ns / 1 ns
module testbench ();
  logic [3:0] s1, s2;
  logic nreset;
  logic lSegEn, rSegEn;
  logic [6:0] seg;
  logic [4:0] sum;
  lab2_vk #('d2) dut (
      .s1(s1),
      .s2(s2),
      .nreset(nreset),
      .lSegEn(lSegEn),
      .rSegEn(rSegEn),
      .seg(seg),
      .sum(sum)
  );

  logic clk;
  assign clk = dut.clk;

  logic lSegEn;
  assign lSegEn = dut.lSegEn;
  logic oldlSegEn;

  int testCounter;
  int errors;

  logic lSegEnExpected;
  logic rSegEnExpected;
  logic [6:0] segExpected;
  logic [4:0] sumExpected;
  logic [21:0] testVectors[1000:0];


  initial begin
    $display("reading test vectors");
    $readmemb("testbench.tv", testVectors);
    testCounter = 0;
    errors = 0;
    nreset = 0;
    #27;
    oldlSegEn = lSegEn;
    nreset = 1;
    #2;
  end

  always @(posedge clk) begin
    #1;
    if (oldlSegEn !== lSegEn) begin
      {s1, s2, lSegEnExpected, rSegEnExpected, segExpected, sumExpected} = testVectors[testCounter];
    end
  end

  always @(negedge clk) begin
    #1;
    if (oldlSegEn !== lSegEn) begin
      if ({lSegEn, rSegEn, seg, sum} !== {lSegEnExpected, rSegEnExpected, segExpected, sumExpected}) begin
        $display("Error (test %d): inputs = %b, %b ", errors, s1, s2);
        $display(
            "outputs = %b segment; L: %b R: %b; %b sum. Expected: (%b segment; L: %b R: %b; %b sum)",
            seg, lSegEn, rSegEn, sum, segExpected, lSegEnExpected, rSegEnExpected, sumExpected);
        errors = errors + 1;
      end
      oldlSegEn   = lSegEn;
      testCounter = testCounter + 1;
      if (testVectors[testCounter] === 22'bx) begin
        $display("%d tests completed with %d errors", testCounter, errors);
        $finish;
      end
    end
  end
endmodule
